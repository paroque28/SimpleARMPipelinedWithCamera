localparam  IMG_WIDTH		=	200;
localparam	IMG_HEIGHT		=	200;
localparam	IMG_PIXELS		=	IMG_WIDTH*IMG_HEIGHT;
localparam  PIXELS          =   $clog2(IMG_HEIGHT*IMG_WIDTH);
