module pipeReg(
	input logic clk,
	input logic rst,
	input logic 
)