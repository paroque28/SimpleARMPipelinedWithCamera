parameter fADD	     = 4'b0000;
parameter fSUB	     = 4'b0001;
parameter fMULT	     = 4'b0010;
parameter fLOAD	     = 4'b0100;
parameter fSTR	     = 4'b0101;
parameter fSL	     = 4'b0110;
parameter fSR	     = 4'b0111;
parameter fB	     = 4'b1000;
parameter fPIC	     = 4'b1001;
parameter fAVERAGE	 = 4'b1010;
parameter fLDA	     = 4'b1011;
parameter fSTR_ONE   = 4'b1100;
parameter fTHI       = 4'b1100;
