localparam  IMG_WIDTH		=	320;
localparam	IMG_HEIGHT		=	240;
localparam	IMG_PIXELS		=	IMG_WIDTH*IMG_HEIGHT;
localparam  PIXELS          =   $clog2(IMG_HEIGHT*IMG_WIDTH);
