parameter BUFFER = 4'b0000;
parameter ADD	 = 4'b0001;
parameter SUB   = 4'b0010;
parameter MULT   = 4'b0011;
parameter DIV	 = 4'b0100;
parameter SL     = 4'b0101;
parameter SR     = 4'b0110;
parameter AV     = 4'b0111;
parameter THI    = 4'b1000;
parameter AND	 = 4'b1001;
parameter NOP	 = 4'b1010;
parameter ORR	 = 4'b1011;
