module pipeReg(
	input logic clk,
	input logic rst,
	input logic enable,
	input logic dataIn[0:31],
	output logic dataOut[0:31]
	
);

endmodule 