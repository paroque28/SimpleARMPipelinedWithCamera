// video.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module video (
		output wire  lcd_clk_clk,        //      lcd_clk.clk
		input  wire  ref_clk_clk,        //      ref_clk.clk
		input  wire  ref_reset_reset,    //    ref_reset.reset
		output wire  reset_source_reset, // reset_source.reset
		output wire  video_in_clk_clk    // video_in_clk.clk
	);

	video_video_pll_0 video_pll_0 (
		.ref_clk_clk        (ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),    //    ref_reset.reset
		.video_in_clk_clk   (video_in_clk_clk),   // video_in_clk.clk
		.lcd_clk_clk        (lcd_clk_clk),        //      lcd_clk.clk
		.reset_source_reset (reset_source_reset)  // reset_source.reset
	);

endmodule
