module memory ();
endmodule 