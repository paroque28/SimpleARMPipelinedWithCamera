
module video (
	lcd_clk_clk,
	ref_clk_clk,
	ref_reset_reset,
	reset_source_reset,
	video_in_clk_clk);	

	output		lcd_clk_clk;
	input		ref_clk_clk;
	input		ref_reset_reset;
	output		reset_source_reset;
	output		video_in_clk_clk;
endmodule
