module memory ()
