localparam FNOP	    = 4'b0000;
localparam FMULT	    = 4'b0001;
localparam FSUB	    = 4'b0010;
localparam FLOAD	    = 4'b0011;
localparam FADD	    = 4'b0100;
localparam FSTR	    = 4'b0101;
localparam FSL	       = 4'b0110;
localparam FSR	       = 4'b0111;
localparam FB	       = 4'b1000;
localparam FPIC	    = 4'b1001;
localparam FAVERAGE	 = 4'b1010;
localparam FLDA	    = 4'b1011;
localparam FORR	    = 4'b1100;
localparam FSTR_ONE   = 4'b1101;
localparam FTHI       = 4'b1111;


localparam OPDATA       = 2'b00;
localparam OPMEMORY     = 2'b01;
localparam OPBRANCH     = 2'b10;
