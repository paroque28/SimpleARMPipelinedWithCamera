module Control_unit (input logic [3:0] opcode,
							
							output logic ALUSrcE,
							output logic [3:0]ALUControlE,
							output logic TfuWD,
							output logic TFUAdd,
							output logic [1:0] MemRd,
							output logic [1:0] MemtoRegW,
							output logic RegSrcD,
							output logic 

							);
							
